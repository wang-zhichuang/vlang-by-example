module main
import hello

fn main() {
	hello.say_hi()
}
